module cpu(clk, reset, s, load, in, out, Z, N, V, w);

endmodule